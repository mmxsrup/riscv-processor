package src_b_mux_pkg;

	localparam SEL_SRC_B_WIDTH = 3;

	localparam SEL_SRC_B_RS2 = 3'h1;
	localparam SEL_SRC_B_IMM = 3'h2;
	localparam SEL_SRC_B_0 = 3'h3;
	localparam SEL_SRC_B_4 = 3'h4;
	localparam SEL_SRC_B_NONE = 3'h0;

endpackage
