package src_a_mux_pkg;

	localparam SEL_SRC_A_WIDTH = 2;

	localparam SEL_SRC_A_PC  = 2'h1;
	localparam SEL_SRC_A_RS1 = 2'h2;
	localparam SEL_SRC_A_IMM = 2'h3;
	localparam SEL_SRC_A_NONE = 2'h0;

endpackage
