package ram_pkg;

	localparam AWIDTH = 32;
	localparam DWIDTH = 32;
	localparam LWIDTH = 4;

endpackage
